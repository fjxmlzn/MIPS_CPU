`timescale 1ns/1ps

module ROM (addr,data);
	input [31:0] addr;
	output [31:0] data;
	reg [31:0] data;
	localparam ROM_SIZE = 32;
	reg [31:0] ROM_DATA[ROM_SIZE-1:0];

	always@(*)
		case(addr[9:2])	//Address Must Be Word Aligned.
			8'd0: data = 32'h08000087;	// j	 entry_main
			8'd1: data = 32'h08000005;	// j	 timer_interrupt_main
			8'd2: data = 32'h0800005e;	// j	 exception_main
			8'd3: data = 32'h08000063;	// j	 uart_send_interrupt_main
			8'd4: data = 32'h08000067;	// j	 uart_recv_interrupt_main
			8'd5: data = 32'h3c084000;	// lui	 $t0, 0x4000
			8'd6: data = 32'h21080008;	// addi	 $t0, $t0, 0x0008
			8'd7: data = 32'h8d090000;	// lw	 $t1, 0, $t0
			8'd8: data = 32'h3129fff9;	// andi	 $t1, $t1, 0xfff9
			8'd9: data = 32'had090000;	// sw	 $t1, 0, $t0
			8'd10: data = 32'h200f00fc;	// addi	 $t7, $zero, 0x00fc
			8'd11: data = 32'h8dea0000;	// lw	 $t2, 0, $t7
			8'd12: data = 32'h8d0b000c;	// lw	 $t3, 12, $t0
			8'd13: data = 32'h000b5a02;	// srl	 $t3, $t3, 8
			8'd14: data = 32'h316c0001;	// andi	 $t4, $t3, 0x0001
			8'd15: data = 32'h000c60c0;	// sll	 $t4, $t4, 3
			8'd16: data = 32'h000b5842;	// srl	 $t3, $t3, 1
			8'd17: data = 32'h016c5825;	// or	 $t3, $t3, $t4
			8'd18: data = 32'h01606020;	// add	 $t4, $t3, $zero
			8'd19: data = 32'h318d0008;	// andi	 $t5, $t4, 0x0008
			8'd20: data = 32'h11a00004;	// beq	 $t5, $zero, ti_getnum
			8'd21: data = 32'h000d6842;	// srl	 $t5, $t5, 1
			8'd22: data = 32'h000a5102;	// srl	 $t2, $t2, 4
			8'd23: data = 32'h01ac6824;	// and	 $t5, $t5, $t4
			8'd24: data = 32'h08000014;	// j	 ti_right_shift_loop
			8'd25: data = 32'h314a000f;	// andi	 $t2, $t2, 0x000f
			8'd26: data = 32'h000b5a00;	// sll	 $t3, $t3, 8
			8'd27: data = 32'h200e0000;	// addi	 $t6, $zero, 0x0
			8'd28: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n0
			8'd29: data = 32'h200e0001;	// addi	 $t6, $zero, 0x1
			8'd30: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n1
			8'd31: data = 32'h200e0002;	// addi	 $t6, $zero, 0x2
			8'd32: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n2
			8'd33: data = 32'h200e0003;	// addi	 $t6, $zero, 0x3
			8'd34: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n3
			8'd35: data = 32'h200e0004;	// addi	 $t6, $zero, 0x4
			8'd36: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n4
			8'd37: data = 32'h200e0005;	// addi	 $t6, $zero, 0x5
			8'd38: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n5
			8'd39: data = 32'h200e0006;	// addi	 $t6, $zero, 0x6
			8'd40: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n6
			8'd41: data = 32'h200e0007;	// addi	 $t6, $zero, 0x7
			8'd42: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n7
			8'd43: data = 32'h200e0008;	// addi	 $t6, $zero, 0x8
			8'd44: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n8
			8'd45: data = 32'h200e0009;	// addi	 $t6, $zero, 0x9
			8'd46: data = 32'h114e001d;	// beq	 $t2, $t6, ti_n9
			8'd47: data = 32'h200e000a;	// addi	 $t6, $zero, 0xa
			8'd48: data = 32'h114e001d;	// beq	 $t2, $t6, ti_na
			8'd49: data = 32'h200e000b;	// addi	 $t6, $zero, 0xb
			8'd50: data = 32'h114e001d;	// beq	 $t2, $t6, ti_nb
			8'd51: data = 32'h200e000c;	// addi	 $t6, $zero, 0xc
			8'd52: data = 32'h114e001d;	// beq	 $t2, $t6, ti_nc
			8'd53: data = 32'h200e000d;	// addi	 $t6, $zero, 0xd
			8'd54: data = 32'h114e001d;	// beq	 $t2, $t6, ti_nd
			8'd55: data = 32'h200e000e;	// addi	 $t6, $zero, 0xe
			8'd56: data = 32'h114e001d;	// beq	 $t2, $t6, ti_ne
			8'd57: data = 32'h08000058;	// j	 ti_nf
			8'd58: data = 32'h216b00fc;	// addi	 $t3, $t3, 0x00fc
			8'd59: data = 32'h0800005a;	// j	 ti_display
			8'd60: data = 32'h216b0060;	// addi	 $t3, $t3, 0x0060
			8'd61: data = 32'h0800005a;	// j	 ti_display
			8'd62: data = 32'h216b00da;	// addi	 $t3, $t3, 0x00da
			8'd63: data = 32'h0800005a;	// j	 ti_display
			8'd64: data = 32'h216b00f2;	// addi	 $t3, $t3, 0x00f2
			8'd65: data = 32'h0800005a;	// j	 ti_display
			8'd66: data = 32'h216b0066;	// addi	 $t3, $t3, 0x0066
			8'd67: data = 32'h0800005a;	// j	 ti_display
			8'd68: data = 32'h216b00b6;	// addi	 $t3, $t3, 0x00b6
			8'd69: data = 32'h0800005a;	// j	 ti_display
			8'd70: data = 32'h216b00be;	// addi	 $t3, $t3, 0x00be
			8'd71: data = 32'h0800005a;	// j	 ti_display
			8'd72: data = 32'h216b00e0;	// addi	 $t3, $t3, 0x00e0
			8'd73: data = 32'h0800005a;	// j	 ti_display
			8'd74: data = 32'h216b00fe;	// addi	 $t3, $t3, 0x00fe
			8'd75: data = 32'h0800005a;	// j	 ti_display
			8'd76: data = 32'h216b00f6;	// addi	 $t3, $t3, 0x00f6
			8'd77: data = 32'h0800005a;	// j	 ti_display
			8'd78: data = 32'h216b00ee;	// addi	 $t3, $t3, 0x00ee
			8'd79: data = 32'h0800005a;	// j	 ti_display
			8'd80: data = 32'h216b00ff;	// addi	 $t3, $t3, 0x00ff
			8'd81: data = 32'h0800005a;	// j	 ti_display
			8'd82: data = 32'h216b009c;	// addi	 $t3, $t3, 0x009c
			8'd83: data = 32'h0800005a;	// j	 ti_display
			8'd84: data = 32'h216b00fd;	// addi	 $t3, $t3, 0x00fd
			8'd85: data = 32'h0800005a;	// j	 ti_display
			8'd86: data = 32'h216b009e;	// addi	 $t3, $t3, 0x009e
			8'd87: data = 32'h0800005a;	// j	 ti_display
			8'd88: data = 32'h216b008e;	// addi	 $t3, $t3, 0x008e
			8'd89: data = 32'h0800005a;	// j	 ti_display
			8'd90: data = 32'had0b000c;	// sw	 $t3, 12, $t0
			8'd91: data = 32'h21290002;	// addi	 $t1, $t1, 2
			8'd92: data = 32'had090000;	// sw	 $t1, 0, $t0
			8'd93: data = 32'h03400008;	// jr	 $26
			8'd94: data = 32'h3c084000;	// lui	 $t0, 0x4000
			8'd95: data = 32'h21080018;	// addi	 $t0, $t0, 0x0018
			8'd96: data = 32'h2009005a;	// addi	 $t1, $zero, 0x005a
			8'd97: data = 32'had090000;	// sw	 $t1, 0, $t0
			8'd98: data = 32'h03400008;	// jr	 $26
			8'd99: data = 32'h3c084000;	// lui	 $t0, 0x4000
			8'd100: data = 32'h21080018;	// addi	 $t0, $t0, 0x0018
			8'd101: data = 32'h8d090000;	// lw	 $t1, 0, $t0
			8'd102: data = 32'h03400008;	// jr	 $26
			8'd103: data = 32'h3c084000;	// lui	 $t0, 0x4000
			8'd104: data = 32'h2108001c;	// addi	 $t0, $t0, 0x001c
			8'd105: data = 32'h8d090000;	// lw	 $t1, 0, $t0
			8'd106: data = 32'h200a00fc;	// addi	 $t2, $zero, 0x00fc
			8'd107: data = 32'h8d4b0000;	// lw	 $t3, 0, $t2
			8'd108: data = 32'h000b6402;	// srl	 $t4, $t3, 16
			8'd109: data = 32'h15800004;	// bne	 $t4, $zero, ur_gcd_start
			8'd110: data = 32'h3c0b0001;	// lui	 $t3, 0x0001
			8'd111: data = 32'h01695820;	// add	 $t3, $t3, $t1
			8'd112: data = 32'had4b0000;	// sw	 $t3, 0, $t2
			8'd113: data = 32'h03400008;	// jr	 $26
			8'd114: data = 32'h00094a00;	// sll	 $t1, $t1, 8
			8'd115: data = 32'h01695820;	// add	 $t3, $t3, $t1
			8'd116: data = 32'h000b5c00;	// sll	 $t3, $t3, 16
			8'd117: data = 32'h000b5c02;	// srl	 $t3, $t3, 16
			8'd118: data = 32'had4b0000;	// sw	 $t3, 0, $t2
			8'd119: data = 32'h316e00ff;	// andi	 $t6, $t3, 0x00ff
			8'd120: data = 32'h316fff00;	// andi	 $t7, $t3, 0xff00
			8'd121: data = 32'h000f7a02;	// srl	 $t7, $t7, 8
			8'd122: data = 32'h11e00007;	// beq	 $t7, $zero, ur_gcd_end
			8'd123: data = 32'h01ee6822;	// sub	 $t5, $t7, $t6
			8'd124: data = 32'h1da00001;	// bgtz	 $t5, ur_gcd_main_swap
			8'd125: data = 32'h01cf7022;	// sub	 $t6, $t6, $t7
			8'd126: data = 32'h000e6820;	// add	 $t5, $zero, $t6
			8'd127: data = 32'h000f7020;	// add	 $t6, $zero, $t7
			8'd128: data = 32'h000d7820;	// add	 $t7, $zero, $t5
			8'd129: data = 32'h0800007a;	// j	 ur_gcd_main
			8'd130: data = 32'h3c084000;	// lui	 $t0, 0x4000
			8'd131: data = 32'h2108000c;	// addi	 $t0, $t0, 0x000c
			8'd132: data = 32'had0e0000;	// sw	 $t6, 0, $t0
			8'd133: data = 32'had0e000c;	// sw	 $t6, 12, $t0
			8'd134: data = 32'h03400008;	// jr	 $26
			8'd135: data = 32'h3c084000;	// lui	 $t0, 0x4000
			8'd136: data = 32'h200907ff;	// addi	 $t1, $zero, 0x07ff
			8'd137: data = 32'had090014;	// sw	 $t1, 0x14, $t0
			8'd138: data = 32'had00000c;	// sw	 $zero, 0x0c, $t0
			8'd139: data = 32'h3c09fffe;	// lui	 $t1, 0xfffe
			8'd140: data = 32'h2129795f;	// addi	 $t1, $t1, 0x795f
			8'd141: data = 32'had090000;	// sw	 $t1, 0, $t0
			8'd142: data = 32'h00004827;	// nor	 $t1, $0, $0
			8'd143: data = 32'had090004;	// sw	 $t1, 0x04, $t0
			8'd144: data = 32'h20090003;	// addi	 $t1, $zero, 0x0003
			8'd145: data = 32'had090008;	// sw	 $t1, 0x08, $t0
			8'd146: data = 32'h20090002;	// addi	 $t1, $zero, 0x0002
			8'd147: data = 32'had090020;	// sw	 $t1, 0x20, $t0
			8'd148: data = 32'h200a0258;	// addi	 $t2, $zero, 0x0254
			8'd149: data = 32'h01400008;	// jr	 $t2
			8'd150: data = 32'hfac23e4e;
			8'd151: data = 32'h08000097;	// j	 main_loop
			default:	data = 32'h08000097;
		endcase
endmodule
